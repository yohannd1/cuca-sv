module tb_ram;
  // TODO

  initial begin
    $display("omg");
    $finish;
  end
endmodule

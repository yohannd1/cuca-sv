module register(
  input logic clock, enable, rw,
  inout logic[BITW-1:0] bus
);

endmodule;

module tb_ram;
  // TODO
endmodule

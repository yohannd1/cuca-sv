module param;
endmodule
